`default_nettype none

module mmu_feeder (
    input wire clk,
    input wire rst,
    input wire en,
    input wire [2:0] mmu_cycle,

    input wire transpose,

    /* Memory module interface */
    input wire [7:0] weight0, weight1, weight2, weight3,
    input wire [7:0] input0, input1, input2, input3,

    /* systolic array -> feeder */
    input wire signed [11:0] c00, c01, c10, c11,

    /* feeder -> mmu */
    output wire clear,
    output reg [7:0] a_data0,
    output reg [7:0] a_data1,
    output reg [7:0] b_data0,
    output reg [7:0] b_data1,

    /* feeder -> rpi */
    output wire done,
    output reg [7:0] host_outdata
);

    // Done signal for output phase
    assign done = en && (mmu_cycle >= 3'b010) && (mmu_cycle <= 3'b101);
    assign clear = (mmu_cycle == 3'b110);

    // Output counter for selecting c_out
    reg [1:0] output_count;

    function [7:0] saturate_to_s8;
        input signed [11:0] val;
        begin
            if (val > 127)
                saturate_to_s8 = 8'sd127;
            else if (val < -128)
                saturate_to_s8 = -8'sd128;
            else
                saturate_to_s8 = val[7:0];
        end
    endfunction

    // Sequential logic for control and data outputs
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            a_data0 <= 0;
            a_data1 <= 0;
            b_data0 <= 0;
            b_data1 <= 0;
            output_count <= 0;
        end else begin
            output_count <= 0;
            if (en) begin
                $display("mmu cycle %d, output count %d", mmu_cycle, output_count);
                $display("a_data0 %d, a_data1 %d, b_data0 %d, b_data1 %d", a_data0, a_data1, b_data0, b_data1);
                // Update output_count during output phase
                if (mmu_cycle >= 3) begin
                    output_count <= output_count + 1;
                end else begin
                    output_count <= 0;
                end
                case (mmu_cycle)
                    3'b000: begin
                        a_data0 <= weight0;
                        b_data0 <= input0;
                    end
                    3'b001: begin
                        a_data0 <= weight1;
                        a_data1 <= weight2;
                        if (transpose) begin
                            b_data0 <= input1;
                            b_data1 <= input2;
                        end else begin
                            b_data0 <= input2;
                            b_data1 <= input1;
                        end
                    end
                    3'b010: begin
                        a_data0 <= 0;
                        a_data1 <= 0;
                        b_data0 <= 0;
                        b_data1 <= input3;
                    end
                    3'b011: begin
                        a_data0 <= 0;
                        b_data1 <= input3;
                        b_data0 <= 0;
                        a_data1 <= weight3;
                    end
                    3'b100: begin
                        a_data0 <= 0;
                        b_data1 <= input3;
                        b_data0 <= 0;
                        a_data1 <= a_data1;
                    end
                    // Other cycles (3'b100 to 3'b101) keep defaults (0)
                    default: begin 
                        a_data0 <= 0;
                        a_data1 <= 0;
                        b_data0 <= 0;
                        b_data1 <= 0;
                    end
                endcase
            end else begin
                a_data0 <= 0;
                a_data1 <= 0;
                b_data0 <= 0;
                b_data1 <= 0;
            end
        end
    end

    // Combinational logic for host_outdata with corrected saturation
    always @(*) begin
        host_outdata = 8'b0; // Default to avoid latch
        if (en) begin
            case (output_count)
                2'b00: host_outdata = saturate_to_s8(c00);
                2'b01: host_outdata = saturate_to_s8(c01);
                2'b10: host_outdata = saturate_to_s8(c10);
                2'b11: host_outdata = saturate_to_s8(c11);
                default: host_outdata = 8'b0;
            endcase
        end
    end

endmodule