module buffer (
    input wire A,
    output wire X
);
    assign X = A;
endmodule